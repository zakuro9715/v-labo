module mod

pub enum Enum {
	value
}

pub fn f(v Enum) {
	println(v)
}
